*---------- DMTH4005SK3 Spice Model ----------
.SUBCKT DMTH4005SK3 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 NMOS L = 1E-006 W = 1E-006 
RD 10 1 9.814E-005 
RS 30 3 0.001 
RG 20 2 0.67 
CGS 2 3 2.961E-009 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1 VFB 1 
CGD 13 14 1.3E-009 
R1 13 0 1 
D1 12 13 DLIM 
DDG 15 14 DCGD 
R2 12 15 1 
D2 15 0 DLIM 
DSD 3 10 DSUB 
.MODEL NMOS NMOS LEVEL = 3 VMAX = 5.378E+005 ETA = 0.001 VTO = 3.117 
+ TOX = 6E-008 NSUB = 1E+016 KP = 46.39 U0 = 400 KAPPA = 10 
.MODEL DCGD D CJO = 1.053E-009 VJ = 0.8 M = 0.6001 
.MODEL DSUB D IS = 1.159E-009 N = 1.284 RS = 0.0003205 BV = 40 CJO = 1.784E-009 VJ = 0.8 M = 0.6 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMTH4005SK3 Spice Model v1.0M Last Revised 2016/3/8