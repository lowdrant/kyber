*SRC=BZT52C2V4LP;BZT52C2V4LP;Diodes;Zener <=10V; 2.40V  0.250W   DIODES ZENER DIODE
*SYM=HZEN
.SUBCKT BZT52C2V4LP  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 0.2
.MODEL DF D ( IS=42.9p RS=35.1 N=1.10
+ CJO=159p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=150n RS=6.5 N=8.0 )
.ENDS