*SRC=BZT52C9V1LP;DI_BZT52C9V1LP;Diodes;Zener <=10V; 9.10V  0.250W   Diodes Inc. QFN Zener
*SYM=HZEN
.SUBCKT DI_BZT52C9V1LP  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 7.44
.MODEL DF D ( IS=11.3p RS=31.3 N=1.10
+ CJO=50.3p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=2.26f RS=3.45 N=2.23 )
.ENDS