*---------- DMP3028LK3 Spice Model ----------
.SUBCKT DMP3028LK3 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 0.01205 
RS 30 3 0.001 
RG 20 2 14.8 
CGS 2 3 1.141E-009 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 8E-010 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 1E-009 
+ TOX = 6E-008 NSUB = 1E+016 KP = 24.29 KAPPA = 55.87 VTO = -2.147 
.MODEL DCGD D CJO = 4.573E-010 VJ = 0.4119 M = 0.3922 
.MODEL DSUB D IS = 2.24E-010 N = 1.262 RS = 0.009108 
+ BV = 50 CJO = 2.261E-010 VJ = 0.5048 M = 0.5435 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMP3028LK3 Spice Model v1.0 Last Revised 2018/2/1